`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/06/2020 12:21:06 PM
// Design Name: 
// Module Name: state_startandgameover
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module state_startandgameover(
        input [9:0] x,
        input [9:0] y,
        output reg tmp
    );
        reg T1;
        reg T2;
    
        reg H1;
        reg H2;
        reg H3;
    
        reg E1;
        reg E2;
        reg E3;
        reg E4;
    
        reg S1;
        reg S2;
        reg S3;
        reg S4;
        reg S5;
        reg S6;
        reg S7;
    
        reg N1;
        reg N2;
        reg N3;
        reg N4;
        reg N5;
        
        reg A1;
        reg A2;
        reg A3;
        reg A4;
    
        reg K1;
        reg K2;
        reg K3;
        reg K4;
        reg K5;
        reg K6;
   
        reg E5;
        reg E6;
        reg E7;
        reg E8;    
        
        reg p1;
        reg p2;
        reg p3;
        reg p4;
        
        reg r1;
        reg r2;
        reg r3;
        reg r4;
        reg r5;
        
        reg ee1;
        reg ee2;
        reg ee3;
        reg ee4;
        
        reg sz1;
        reg sz2;
        reg sz3;
        reg sz4;
        reg sz5;
        reg sz6;
        reg sz7;
        reg sz8;
        reg sz9;
        reg sz10;
        reg sz11;
        reg sz12;
        reg sz13;
        reg sz14;
        
        reg aa1;
        reg aa2;
        reg aa3;
        reg aa4;
        
        reg nn1;
        reg nn2;
        reg nn3;
        reg nn4;
        reg nn5;
        
        reg yy1;
        reg yy2;
        reg yy3;
        reg yy4;
        reg yy5;
        
        reg bb1;
        reg bb2;
        reg bb3;
        reg bb4;
        reg bb5;
        reg bb6;
        
        reg o1;
        reg o2;
        reg o3;
        reg o4;
        
        reg t1;
        reg t2;
        
        reg t3;
        reg t4;
        
        reg o5;
        reg o6;
        reg o7;
        reg o8;
        
        reg nn6;
        reg nn7;
        reg nn8;
        reg nn9;
        reg nn10;
        
        reg t5;
        reg t6;
        
        reg o9;
        reg o10;
        reg o11;
        reg o12;
        
        reg sz15;
        reg sz16;
        reg sz17;
        reg sz18;
        reg sz19;
        reg sz20;
        reg sz21;
        
        reg t7;
        reg t8;
        
        reg aa5;
        reg aa6;
        reg aa7;
        reg aa8;
        
        reg r6;
        reg r7;
        reg r8;
        reg r9;
        reg r10;
        
        reg t9;
        reg t10;
        
    always@(*)
    begin
        //T
        T1 = ((x>125) & (x<=165)) & ((y>120) & (y<=130));
        T2 = ((x>140) & (x<=150)) & ((y>=131) & (y<=200));
        //H
        H1 = ((x>=171) & (x<=180)) & ((y>120) & (y<=200));
        H2 = ((x>=171) & (x<=210)) & ((y>155) & (y<=165));
        H3 = ((x>=201) & (x<=210)) & ((y>120) & (y<=200));
        //E
        E1 = ((x>=216) & (x<=225)) & ((y>=121) & (y<=200));
        E2 = ((x>=226) & (x<=255)) & ((y>=121) & (y<=130));
        E3 = ((x>=226) & (x<=255)) & ((y>=156) & (y<=165));
        E4 = ((x>=226) & (x<=255)) & ((y>=191) & (y<=200));
        //S
        S1 = ((x>=296) & (x<=305)) & ((y>=131) & (y<=155));
        S2 = ((x>=306) & (x<=325)) & ((y>=121) & (y<=130));
        S3 = ((x>=326) & (x<=335)) & ((y>=131) & (y<=143));
        S4 = ((x>=306) & (x<=325)) & ((y>=156) & (y<=165));
        S5 = ((x>=326) & (x<=335)) & ((y>=166) & (y<=190));
        S6 = ((x>=306) & (x<=325)) & ((y>=191) & (y<=200));
        S7 = ((x>=296) & (x<=305)) & ((y>=178) & (y<=190));
        //N
        N1 = ((x>=341) & (x<=348)) & ((y>=121) & (y<=200));
        N2 = ((x>=349) & (x<=356)) & ((y>=131) & (y<=151));
        N3 = ((x>=357) & (x<=364)) & ((y>=156) & (y<=165));
        N4 = ((x>=365) & (x<=372)) & ((y>=166) & (y<=190));
        N5 = ((x>=373) & (x<=380)) & ((y>=121) & (y<=200));
        //A
        A1 = ((x>=386) & (x<=395)) & ((y>=131) & (y<=200));
        A2 = ((x>=396) & (x<=415)) & ((y>=121) & (y<=130));
        A3 = ((x>=396) & (x<=415)) & ((y>=161) & (y<=170));
        A4 = ((x>=416) & (x<=425)) & ((y>=131) & (y<=200));
        //K
        K1 = ((x>=431) & (x<=440)) & ((y>=121) & (y<=200));
        K2 = ((x>=441) & (x<=450)) & ((y>=156) & (y<=165));
        K3 = ((x>=461) & (x<=470)) & ((y>=121) & (y<=145));
        K4 = ((x>=451) & (x<=460)) & ((y>=146) & (y<=155));
        K5 = ((x>=451) & (x<=460)) & ((y>=166) & (y<=175));
        K6 = ((x>=461) & (x<=470)) & ((y>=176) & (y<=200));
        //E
        E5 = ((x>=476) & (x<=485)) & ((y>=121) & (y<=200));
        E6 = ((x>=486) & (x<=515)) & ((y>=121) & (y<=130));
        E7 = ((x>=486) & (x<=515)) & ((y>=156) & (y<=165));
        E8 = ((x>=486) & (x<=515)) & ((y>=191) & (y<=200));
        
        //P
        p1 = ((x>=46) & (x<=50)) & ((y>=321) & (y<=360));
        p2 = ((x>=51) & (x<=60)) & ((y>=321) & (y<=325));
        p3 = ((x>=51) & (x<=60)) & ((y>=341) & (y<=345));
        p4 = ((x>=61) & (x<=65)) & ((y>=326) & (y<=340));
        //R
        r1 = ((x>=69) & (x<=73)) & ((y>=321) & (y<=360));
        r2 = ((x>=74) & (x<=83)) & ((y>=321) & (y<=325));
        r3 = ((x>=74) & (x<=83)) & ((y>=341) & (y<=345));
        r4 = ((x>=84) & (x<=88)) & ((y>=326) & (y<=340));
        r5 = ((x>=84) & (x<=88)) & ((y>=346) & (y<=360));
        //E
        ee1 = ((x>=92) & (x<=96)) & ((y>=321) & (y<=360));
        ee2 = ((x>=97) & (x<=111)) & ((y>=321) & (y<=325));
        ee3 = ((x>=97) & (x<=111)) & ((y>=338) & (y<=343));
        ee4 = ((x>=97) & (x<=111)) & ((y>=356) & (y<=360));
        //S
        sz1 = ((x>=115) & (x<=119)) & ((y>=326) & (y<=338));
        sz2 = ((x>=120) & (x<=129)) & ((y>=321) & (y<=325));
        sz3 = ((x>=130) & (x<=134)) & ((y>=326) & (y<=329));
        sz4 = ((x>=120) & (x<=129)) & ((y>=339) & (y<=343));
        sz5 = ((x>=130) & (x<=134)) & ((y>=344) & (y<=355));
        sz6 = ((x>=120) & (x<=129)) & ((y>=356) & (y<=360));
        sz7 = ((x>=115) & (x<=119)) & ((y>=352) & (y<=355));
        //S
        sz8 = ((x>=138) & (x<=144)) & ((y>=328) & (y<=337));
        sz9 = ((x>=145) & (x<=150)) & ((y>=321) & (y<=327));
        sz10 = ((x>=151) & (x<=157)) & ((y>=328) & (y<=331));
        sz11 = ((x>=145) & (x<=150)) & ((y>=338) & (y<=343));
        sz12 = ((x>=151) & (x<=157)) & ((y>=344) & (y<=353));
        sz13 = ((x>=145) & (x<=150)) & ((y>=354) & (y<=360));
        sz14 = ((x>=138) & (x<=144)) & ((y>=350) & (y<=353));
        //A
        aa1 = ((x>=178) & (x<=182)) & ((y>=326) & (y<=360));
        aa2 = ((x>=183) & (x<=192)) & ((y>=321) & (y<=325));
        aa3 = ((x>=183) & (x<=192)) & ((y>=339) & (y<=343));
        aa4 = ((x>=193) & (x<=197)) & ((y>=326) & (y<=360));
        //N
        nn1 = ((x>=201) & (x<=204)) & ((y>=321) & (y<=360));
        nn2 = ((x>=205) & (x<=208)) & ((y>=326) & (y<=338));
        nn3 = ((x>=209) & (x<=212)) & ((y>=339) & (y<=343));
        nn4 = ((x>=213) & (x<=216)) & ((y>=344) & (y<=355));
        nn5 = ((x>=217) & (x<=220)) & ((y>=321) & (y<=360));
        //Y
        yy1 = ((x>=224) & (x<=227)) & ((y>=321) & (y<=333));
        yy2 = ((x>=228) & (x<=231)) & ((y>=334) & (y<=345));
        yy3 = ((x>=232) & (x<=235)) & ((y>=346) & (y<=360));
        yy4 = ((x>=236) & (x<=239)) & ((y>=334) & (y<=345));
        yy5 = ((x>=240) & (x<=243)) & ((y>=321) & (y<=333));
        //B
        bb1 = ((x>=264) & (x<=268)) & ((y>=321) & (y<=360));
        bb2 = ((x>=269) & (x<=278)) & ((y>=321) & (y<=325));
        bb3 = ((x>=279) & (x<=283)) & ((y>=326) & (y<=338));
        bb4 = ((x>=279) & (x<=283)) & ((y>=344) & (y<=355));
        bb5 = ((x>=269) & (x<=278)) & ((y>=356) & (y<=360));
        bb6 = ((x>=269) & (x<=278)) & ((y>=339) & (y<=343));
        //U
        o1 = ((x>=287) & (x<=291)) & ((y>=321) & (y<=360));
        //o2 = ((x>=292) & (x<=301)) & ((y>=321) & (y<=325));
        o3 = ((x>=302) & (x<=306)) & ((y>=321) & (y<=360));
        o4 = ((x>=292) & (x<=301)) & ((y>=356) & (y<=360));
        //T
        t1 = ((x>=310) & (x<=329)) & ((y>=321) & (y<=330));
        t2 = ((x>=317) & (x<=321)) & ((y>=331) & (y<=360));
        //T
        t3 = ((x>=333) & (x<=352)) & ((y>=321) & (y<=330));
        t4 = ((x>=340) & (x<=344)) & ((y>=331) & (y<=360));
        //O
        o5 = ((x>=356) & (x<=360)) & ((y>=326) & (y<=355));
        o6 = ((x>=361) & (x<=370)) & ((y>=321) & (y<=325));
        o7 = ((x>=371) & (x<=375)) & ((y>=326) & (y<=355));
        o8 = ((x>=361) & (x<=370)) & ((y>=356) & (y<=360));
        //N
        nn6 = ((x>=379) & (x<=382)) & ((y>=321) & (y<=360));
        nn7 = ((x>=383) & (x<=386)) & ((y>=326) & (y<=338));
        nn8 = ((x>=387) & (x<=390)) & ((y>=339) & (y<=343));
        nn9 = ((x>=391) & (x<=394)) & ((y>=344) & (y<=355));
        nn10 = ((x>=395) & (x<=398)) & ((y>=321) & (y<=360));
        //T
        t5 = ((x>=419) & (x<=438)) & ((y>=321) & (y<=330));
        t6 = ((x>=426) & (x<=430)) & ((y>=331) & (y<=360));
        //O
        o9 = ((x>=442) & (x<=446)) & ((y>=326) & (y<=355));
        o10 = ((x>=447) & (x<=456)) & ((y>=321) & (y<=325));
        o11 = ((x>=457) & (x<=461)) & ((y>=326) & (y<=355));
        o12 = ((x>=447) & (x<=456)) & ((y>=356) & (y<=360));
        //S
        sz15 = ((x>=482) & (x<=486)) & ((y>=326) & (y<=338));
        sz16 = ((x>=487) & (x<=496)) & ((y>=321) & (y<=325));
        sz17 = ((x>=497) & (x<=501)) & ((y>=326) & (y<=329));
        sz18 = ((x>=487) & (x<=496)) & ((y>=339) & (y<=343));
        sz19 = ((x>=497) & (x<=501)) & ((y>=344) & (y<=355));
        sz20 = ((x>=487) & (x<=496)) & ((y>=356) & (y<=360));
        sz21 = ((x>=482) & (x<=486)) & ((y>=352) & (y<=355));
        //T
        t7 = ((x>=505) & (x<=524)) & ((y>=321) & (y<=330));
        t8 = ((x>=512) & (x<=516)) & ((y>=331) & (y<=360));
        //A
        aa5 = ((x>=528) & (x<=532)) & ((y>=326) & (y<=360));
        aa6 = ((x>=533) & (x<=542)) & ((y>=321) & (y<=325));
        aa7 = ((x>=533) & (x<=542)) & ((y>=339) & (y<=343));
        aa8 = ((x>=543) & (x<=547)) & ((y>=326) & (y<=360));
        //R
        r6 = ((x>=551) & (x<=555)) & ((y>=321) & (y<=360));
        r7 = ((x>=556) & (x<=565)) & ((y>=321) & (y<=325));
        r8 = ((x>=556) & (x<=565)) & ((y>=341) & (y<=345));
        r9 = ((x>=566) & (x<=570)) & ((y>=326) & (y<=340));
        r10 = ((x>=566) & (x<=570)) & ((y>=346) & (y<=360));
        //T
        t9 = ((x>=574) & (x<=593)) & ((y>=321) & (y<=330));
        t10 = ((x>=581) & (x<=585)) & ((y>=331) & (y<=360));
        
        
        
        tmp = T1 | T2 | H1 | H2 | H3 | E1 | E2 | E3 | E4 | S1 | S2 | S3 | S4 | S5 | S6 | S7 | N1 | N2 | N3 | N4 | N5 | A1 | A2 | A3 | A4 | K1 | K2 | K3 | K4 | K5 | K6 | E5 | E6 | E7 | E8 | p1 | p2 | p3 | p4 | r1 | r2 | r3 | r4 | r5 | ee1 | ee2 | ee3 | ee4 | sz1 | sz2 | sz3 | sz4 | sz5 | sz6 | sz7 | sz8 | sz9 | sz10 | sz11 | sz12 | sz13 | sz14 | aa1 | aa2 | aa3 | aa4 | nn1 | nn2 | nn3 | nn4 | nn5 | yy1 | yy2 | yy3 | yy4 | yy5 | bb1 | bb2 | bb3 | bb4 | bb5 | bb6 | o1 | o2 | o3 | o4 | t1 | t2 | t3 | t4 | o5 | o6 | o7 | o8 | nn6 | nn7 | nn8 | nn9 | nn10 | t5 | t6 | o9 | o10 | o11 | o12 | sz15 | sz16 | sz17 | sz18 | sz19 | sz20 | sz21 | t7 | t8 | aa5 | aa6 | aa7 | aa8 | r6 | r7 | r8 | r9 | r10 | t9 | t10;
    end
    
endmodule
